module AndGate(
    
);

endmodule