module fft_256(
    input clk,
    input rst_n,
    input inv,
    input valid_in.
    input [15:0] x_re,
    input [15:0] x_im,
    output [15:0] y_re,
    output [15:0] y_im
);