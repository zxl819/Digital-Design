module mux4_1(
    input wire[1:0]d0,d1,d2,d3, // 4 inputs
    input wire[1:0]sel,// 2-bit select
    output wire[1:0] mux_out // 2-bit output
);
    always @(*) begin
        
    end
        


endmodule