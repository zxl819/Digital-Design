module seq_circuit2(
    input C,
    input clk,
    input rst_n,
    output wire Y
);
endmodule