module mux4_12(
    input wire sel,
    input [1:0] d1,d2,d3,d0,
    output reg[1:0] out
);

endmodule