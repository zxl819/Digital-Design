module mux4_12(
    input wire sel,
    input [1:0] d1,d2,d3,d0
);

endmodule