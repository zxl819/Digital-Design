module cache_set(
    input wire clk,
    input wire rst_n,
);
