module main_mod();
endmodule

module sub_mod();