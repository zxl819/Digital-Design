module function_mod(
    input [3:0]a,
);