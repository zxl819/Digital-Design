module Tff_22(
    input wire data,
    input wire clk,
    input wire rst,
    output reg q

);

endmodule