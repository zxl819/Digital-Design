module seq_circuit(
    input A,
    input clk,
    input rst_n,
    output wire Y
);


endmodule