module rom(
    input clk,
);
endmodule