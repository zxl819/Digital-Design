module seq_circuit();