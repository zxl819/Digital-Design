module rom(
    input clk,
    input rst_n,
    input [7:0]addr,
    output [3:0]data
);
endmodule