module generted2(
    
);
endmodule