module Tff_2(
    input wire data,clk,rst,
    output reg q
);


endmodule