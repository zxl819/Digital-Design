module main_mod();
endmodule