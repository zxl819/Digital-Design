module seq_circuit(
    input A,
    input clk,
    input rst_n,
    output wire Y
);

reg r0, r1;
always @(posedge clk or negedge rst_n) begin
    
end
endmodule