module main_mod(
    input clk,
    input rst_n,
    input [7:0]a,
    input [7:0]b,
    input [7:0]c,
    
    output [7:0]d
);

endmodule

module sub_mod(
    input clk,
    input rst_n,
    input [7:0]a,
    input [7:0]b,    
    output [7:0]d

);
endmodule