//异步复位串联T触发器
module Tff_2(
    input wire data,clk,rst,
    output reg q
);
always @(posedge clk or negedge rst)

endmodule