module Rom(
    
);
endmodule