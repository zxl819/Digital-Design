module AndGate(
    //input
    input A,
    input B,
    //output
    output Y

);

assign Y = A & B;

endmodule