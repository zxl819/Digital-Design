module odd_sel(
    input [31:0]d,
    input mod_name instance_name (.*);
);
endmodule
