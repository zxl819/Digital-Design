module rom(
    input clk,
    input rst_n,
    input [7:0]addr,
    output [3:0]data
);

reg [3:0]rom[7:0];
always @(posedge clk or negedge rst_n) begin 
    if(~rst_n)begin
        rom[0] <= 4'd0;
        rom[1] <= 4'd2;
        rom[2] <= 4'd4;
        rom[3] <= 4'd6;
        rom[4] <= 4'd8;
        rom[5] <= 4'd10;
        rom[6] <= 4'd12;
    end
end
endmodule