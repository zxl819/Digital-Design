module cache_set(
    input wire clk,
    input wire rst_n,
    input wire [31:0] addr,
    
);
