module cache_set(
    input wire clk,
);
