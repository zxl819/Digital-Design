module generted2(
    input [7:0]data_in,
    input [7:0]data_out
);

genvar i;

endmodule