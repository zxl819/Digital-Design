module seq_circuit();
endmodule