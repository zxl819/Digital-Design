module butterfly(
    input clk, 
    input rst_n,
    input en,
    input signed [15:0] xp_re,
    input signed [15:0] xp_im,
    input signed [15:0] xq_re,
    input signed [15:0] xq_im,
    input signed [15:0] factor_re,
    input signed [15:0] factor_im,
    output vld,
    output signed [15:0] yp_re,
    output signed [15:0] yp_im,
    output signed [15:0] yq_re,
    output signed [15:0] yq_im
);
reg [3:0] en_r;
    //----------------------------------------------------------------------------
    // 1) 使能信号的流水寄存
    //----------------------------------------------------------------------------

always @(posedge clk or negedge rst_n) begin
    if (rst_n == 1'b0) begin
        en_r <= 0;
    end
    else begin
        en_r <= {en_r[2:0], en};
    end
end
assign vld = en_r[2];

//----------------------------------------------------------------------------
// 2) 第 1 拍：计算 xq 与旋转因子的乘积，并把 xp 做移位对齐
//----------------------------------------------------------------------------


reg signed [31:0] xq_wnr_re0;
reg signed [31:0] xq_wnr_re1;
reg signed [31:0] xq_wnr_im0;
reg signed [31:0] xq_wnr_im1;
reg signed [31:0] xp_re_d;
reg signed [31:0] xp_im_d;

always @(posedge clk or negedge rst_n) begin
    if (rst_n == 1'b0) begin
        xp_re_d <= 0;
        xp_im_d <= 0;
        xq_wnr_re0 <= 0;
        xq_wnr_re1 <= 0;
        xq_wnr_im0 <= 0;
        xq_wnr_im1 <= 0;

    end
    else if(en) begin  //bufferfly algorithm
        xq_wnr_re0 <= xq_re * factor_re; 
        xq_wnr_re1 <= xq_im * factor_im;
        xq_wnr_im0 <= xq_re * factor_im;
        xq_wnr_im1 <= xq_im * factor_re;

        //xp 左移15位
        xp_re_d <= {{4{xp_re[15]}}, xp_re[14:0],13'b0};
        xp_im_d <= {{4{xp_im[15]}}, xp_im[14:0],13'b0};
    end
end
    //----------------------------------------------------------------------------
    // 3) 第 2 拍：蝶形核心加/减(合并乘积)
    //----------------------------------------------------------------------------


reg signed [31:0] xq_wnr_re;
reg signed [31:0] xq_wnr_im;
reg signed [31:0] xp_re_d1;
reg signed [31:0] xp_im_d1; 

always @(posedge clk or negedge rst_n) begin
    if (rst_n == 1'b0) begin
        xq_wnr_re <= 0;
        xq_wnr_im <= 0;
        xp_re_d1 <= 0;
        xp_im_d1 <= 0;
    end
    else if(en_r[0]) begin
        xp_re_d1 <= xp_re_d;
        xp_im_d1 <= xp_im_d;
        xq_wnr_re <= xq_wnr_re0 - xq_wnr_re1;// xq * Wn 的实部
        xq_wnr_im <= xq_wnr_im0 + xq_wnr_im1;// xq * Wn 的虚部
    end
end

    //----------------------------------------------------------------------------
    // 4) 第 3 拍：最终蝶形加减(与 xp 相加/相减)
    //----------------------------------------------------------------------------

reg signed [31:0] yp_re_r;
reg signed [31:0] yp_im_r;
reg signed [31:0] yq_re_r;
reg signed [31:0] yq_im_r;

always @(posedge clk or negedge rst_n) begin
    if (rst_n == 1'b0) begin
        yp_re_r <= 0;
        yp_im_r <= 0;
        yq_re_r <= 0;
        yq_im_r <= 0;
    end
    else if(en_r[1]) begin
        yp_re_r <= xp_re_d1 + xq_wnr_re;
        yp_im_r <= xp_im_d1 + xq_wnr_im;
        yq_re_r <= xp_re_d1 - xq_wnr_re;
        yq_im_r <= xp_im_d1 - xq_wnr_im;
    end
end

    assign yp_re = {yp_re_r[31],yp_re_r[13+15:13]};
    assign yp_im = {yp_im_r[31],yp_im_r[13+15:13]};
    assign yq_re = {yq_re_r[31],yq_re_r[13+15:13]};
    assign yq_im = {yq_im_r[31],yq_im_r[13+15:13]};

endmodule