module mux4_1(

    
);

endmodule